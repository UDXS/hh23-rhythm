module sc_engine(
    input clk,
    input reset,
    input req_stb,

    